`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 17.03.2018 15:01:45
// Design Name: 
// Module Name: nuevo
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

primera prueba

edicion numero 2 Ronny Zarate

edicion número 3 Ronny Zarate

module nuevo(

    );
endmodule
